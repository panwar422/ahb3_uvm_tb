`define COUNT 7

typedef enum bit [1:0] {IDLE, BUSY, NONSEQ, SEQ} transfer_t;
typedef enum bit {READ,WRITE} rw_t;
typedef enum bit [2:0] {SINGLE, INCR, WRAP4, INCR4, WRAP8, INCR8, WRAP16, INCR16} burst_t;
typedef enum bit [2:0] {BYTE, HALFWORD, WORD, WORDx2, WORDx4, WORDx8, WORDx16, WORDx32} size_t;
typedef enum bit [1:0] {OKAY, ERROR, RETRY, SPLIT} response_t;

#addind something into it 
